LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY regn IS
    GENERIC (data_width : INTEGER);
    PORT (
        clr : IN STD_LOGIC;
        clk : IN STD_LOGIC;
        en : IN STD_LOGIC;
        d : IN STD_LOGIC_VECTOR(data_width - 1 DOWNTO 0);
        q : OUT STD_LOGIC_VECTOR(data_width - 1 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE behavior OF regn IS
BEGIN
    PROCESS (clr, clk)
    BEGIN
        IF (clr = '1') THEN
            q <= (OTHERS => '0');
        ELSIF (clk'event AND clk = '1' AND en = '1') THEN
            q <= d;
        END IF;
    END PROCESS;
END;